`timescale 1ns/100ps

module Instr_Mem (
    input wire [31:0] addr,  // programming counter addr (motion that should do)
    output reg [31:0] instr  // instr output
);

    reg [31:0] memory [0:65535]; //64k instr = 128kbyte
    // initial (wouldn't change if u don't want to do more)
    initial begin
// ********************整數運算*********************
// opcode rs rs2 rd imm	
//(R-type)
        memory[0]  = 32'b0000000_00011_00010_000_00001_0110011; // add x1, x2, x3
        memory[1]  = 32'b0100000_00011_00010_000_00001_0110011; // sub x1, x2, x3
        memory[2]  = 32'b0000000_00011_00010_100_00001_0110011; // xor x1, x2, x3
        memory[3]  = 32'b0000000_00011_00010_110_00001_0110011; // or x1, x2, x3
        memory[4]  = 32'b0000000_00011_00010_111_00001_0110011; // and x1, x2, x3
        memory[5]  = 32'b0000000_00011_00010_001_00001_0110011; // sll x1, x2, x3
        memory[6]  = 32'b0000000_00011_00010_101_00001_0110011; // srl x1, x2, x3
        memory[7]  = 32'b0100000_00011_00010_101_00001_0110011; // sra x1, x2, x3
        memory[8]  = 32'b0000000_00011_00010_010_00001_0110011; // slt x1, x2, x3
        memory[9]  = 32'b0000000_00011_00010_011_00001_0110011; // sltu x1, x2, x3
        
//(I-type)						       								
        memory[10] = 32'b000000000001_00010_000_00001_0010011; // addi x1, x2, 1
        memory[11] = 32'b000000000001_00010_100_00001_0010011; // xori x1, x2, 1
        memory[12] = 32'b000000000001_00010_110_00001_0010011; // ori x1, x2, 1
        memory[13] = 32'b000000000001_00010_111_00001_0010011; // andi x1, x2, 1
        memory[14] = 32'b000000000001_00010_001_00001_0010011; // slli x1, x2, 1 (shamt) 
        memory[15] = 32'b000000000001_00010_101_00001_0010011; // srli x1, x2, 1 (shamt)
        memory[16] = 32'b010000000001_00010_101_00001_0010011; // srai x1, x2, 1 (shamt)
        memory[17] = 32'b000000000001_00010_010_00001_0010011; // slti x1, x2, 1
        memory[18] = 32'b000000000001_00010_011_00001_0010011; // sltiu x1, x2, 1
//(U-type)
	memory[19] = 32'b000000000001_00010_000_00001_0110111; // lui imm rd 1
        memory[20] = 32'b000000000001_00010_100_00001_0010111; // auipe 
// ********************條件跳轉*********************
// (B-type)
        memory[21] = 32'b0000000_00010_00001_000_00010_1100011; // beq x1, x2, offset
        memory[22] = 32'b0000000_00010_00001_001_00010_1100011; // bne x1, x2, offset
        memory[23] = 32'b0000000_00010_00001_100_00010_1100011; // blt x1, x2, offset
        memory[24] = 32'b0000000_00010_00001_101_00010_1100011; // bge x1, x2, offset
        memory[25] = 32'b0000000_00010_00001_110_00010_1100011; // bltu x1, x2, offset
        memory[26] = 32'b0000000_00010_00001_111_00010_1100011; // bgeu x1, x2, offset
// (J-type)
        memory[27] = 32'b000000000100_00000_110_00001_1101111; // jal x1, offset
        memory[28] = 32'b000000000100_00001_000_00010_1100111; // jalr x2, x1, offset

// ********************reading instru*********************
        memory[29] = 32'b000000000000_00101_010_00100_0000011;  // lw x4, 0(x5)
        memory[30] = 32'b000000000000_00101_000_00100_0000011;  // lb x4, 0(x5)
        memory[31] = 32'b000000000000_00101_001_00100_0000011;  // lh x4, 0(x5)
        memory[32] = 32'b000000000000_00101_100_00100_0000011;  // lbu x4, 0(x5)
        memory[33] = 32'b000000000000_00101_101_00100_0000011;  // lhu x4, 0(x5)
        memory[34] = 32'b0000000_00001_00010_010_00000_0100011; // sw x1, 0(x2)
        memory[35] = 32'b0000000_00001_00010_000_00000_0100011; // sb x1, 0(x2)
        memory[36] = 32'b0000000_00001_00010_001_00000_0100011; // sh x1, 0(x2)

//********************pesudo instr*********************
        memory[37] = 32'b000000000000_00000_000_00000_0010011; // nop (addi x0, x0, 0)
        memory[38] = 32'b000000000000_00001_000_00010_0110011; // mv x2, x1 (add x2, x1, x0)
        memory[39] = 32'b000000000000_00000_000_00001_0010011; // li x1, 0 (addi x1, x0, 0)
        memory[40] = 32'b000000000100_00000_110_00001_1101111; // call (jal x1, offset)
        memory[41] = 32'b000000000000_00001_000_00010_1100111; // ret (jalr x0, x1, 0)


    end
// 共41條指令
    // IF
    always @(*) begin
        instr = memory[addr[17:2]]; // addr[17:2]
	// 2^16 = 65535 
	// 每條指令間隔4bytes +4 > 省略01 ＝ 1 / 00 ＝ 0 / 11 ＝ 3 / 10 ＝ 2 的可能
    end
endmodule

